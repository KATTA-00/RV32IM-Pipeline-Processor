module control()