

module decode_stage_tb;

    


endmodule